** Profile: "SCHEMATIC1-OSC"  [ X:\Projects\Engineering\ProjectScience\hardware\pspice\osc\OSC-PSpiceFiles\SCHEMATIC1\OSC.sim ] 

** Creating circuit file "OSC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\InnovusSollertia\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.STEP LIN V_V1 1 5 0.1 
.TEMP 27
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
